// simple_module.v
module simple_module(input a, input b, output y);
    assign y = a & b;  // AND gate
endmodule

